module cpu(
	input wire [3:0] in,
	input wire clock,
	input wire ZF,
	input wire CF,
	output wire HLT,
	output wire MI,
	output wire RI,
	output wire RO,
	output wire IO,
	output wire II,
	output wire AI,
	output wire AO,
	output wire EO,
	output wire SU,
	output wire BI,
	output wire BO,
	output wire OI,
	output wire CE,
	output wire CO,
	output wire J,
	output wire FI,
	output wire [7:0] BRUH
);

wire [3:0] count_cpu;

assign BO = 0;

counter counter(
	.in(),
	.clock(clock),
	.reset(count_cpu === 6 | reset),
	.jump(),
	.enable(1'b1),
	.out(count_cpu)
);

// Markers for cpu_gen.py, DO NOT DELETE
// START
// Generated by cpu_gen.py at 2021-05-12 22:15:53.312897
// by Jonathan Gai
reg [15:0] out;

assign {HLT, MI, RI, RO, IO, II, AI, AO, EO, SU, BI,
		OI, CE, CO, J, FI} = out;
always @(posedge clock) begin
	case ({in, count_cpu})
		// NOP
		8'b00000000: out <= 16'b0100000000000100;
		8'b00000001: out <= 16'b0001010000001000;
		// LDA
		8'b00010000: out <= 16'b0100000000000100;
		8'b00010001: out <= 16'b0001010000001000;
		8'b00010010: out <= 16'b0100100000000000;
		8'b00010011: out <= 16'b0001001000000000;
		// ADD
		8'b00100000: out <= 16'b0100000000000100;
		8'b00100001: out <= 16'b0001010000001000;
		8'b00100010: out <= 16'b0100100000000000;
		8'b00100011: out <= 16'b0001000000100000;
		8'b00100100: out <= 16'b0000001010000000;
		// SUB
		8'b00110000: out <= 16'b0100000000000100;
		8'b00110001: out <= 16'b0001010000001000;
		8'b00110010: out <= 16'b0100100000000000;
		8'b00110011: out <= 16'b0001000000100000;
		8'b00110100: out <= 16'b0000001011000000;
		// STA
		8'b01000000: out <= 16'b0100000000000100;
		8'b01000001: out <= 16'b0001010000001000;
		8'b01000010: out <= 16'b0100100000000000;
		8'b01000011: out <= 16'b0010000100000000;
		// LDI
		8'b01010000: out <= 16'b0100000000000100;
		8'b01010001: out <= 16'b0001010000001000;
		8'b01010010: out <= 16'b0000101000000000;
		// JMP
		8'b01100000: out <= 16'b0100000000000100;
		8'b01100001: out <= 16'b0001010000001000;
		8'b01100010: out <= 16'b0000100000000010;
		// OUT
		8'b11100000: out <= 16'b0100000000000100;
		8'b11100001: out <= 16'b0001010000001000;
		8'b11100010: out <= 16'b0000000100010000;
		// HLT
		8'b11110000: out <= 16'b0100000000000100;
		8'b11110001: out <= 16'b0001010000001000;
		8'b11110010: out <= 16'b1000000000000000;
		default:     out <= 16'b0000000000000000;
	endcase
end
// FINISH
endmodule
